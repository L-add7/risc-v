`define RF_PATH   riscv.rf
`define DMEM_PATH riscv.dmem
`define IMEM_PATH riscv.imem
